`timescale 1ns/1ps
module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];
always@(*)
	case(addr[10:2])
		0: data <= 32'h08000003;
		1: data <= 32'h08000003;
		2: data <= 32'h08000003;
		3: data <= 32'h200e0024;
		4: data <= 32'h3c024000;
		5: data <= 32'hac400008;
		6: data <= 32'h2004fc18;
		7: data <= 32'hac440000;
		8: data <= 32'h01c00008;
		9: data <= 32'h2004ffff;
		10: data <= 32'hac440004;
		11: data <= 32'h20050003;
		12: data <= 32'hac450008;
		13: data <= 32'h20180008;
		14: data <= 32'h8c430018;
		15: data <= 32'h2063ffff;
		16: data <= 32'h1860fffd;
		17: data <= 32'h8c48001c;
		18: data <= 32'h8c50001c;
		19: data <= 32'h8c490020;
		20: data <= 32'h8c510020;
		21: data <= 32'h01005020;
		22: data <= 32'h01495022;
		23: data <= 32'h1d40fffe;
		24: data <= 32'h11400004;
		25: data <= 32'h01495020;
		26: data <= 32'h01204020;
		27: data <= 32'h01404820;
		28: data <= 32'h08000015;
		29: data <= 32'hac490024;
		30: data <= 32'hac49000c;
		31: data <= 32'h00802020;
		32: data <= 32'h0800001f;
		33: data <= 32'h8c4b0008;
		34: data <= 32'h316bfff9;
		35: data <= 32'hac4b0008;
		36: data <= 32'h20190008;
		37: data <= 32'h1319000d;
		38: data <= 32'h0019c842;
		39: data <= 32'h13190008;
		40: data <= 32'h0019c842;
		41: data <= 32'h13190002;
		42: data <= 32'h0019c842;
		43: data <= 32'h1319000b;
		44: data <= 32'h0010a700;
		45: data <= 32'h0014a702;
		46: data <= 32'h0018c240;
		47: data <= 32'h08000043;
		48: data <= 32'h0010a102;
		49: data <= 32'h0018c240;
		50: data <= 32'h08000043;
		51: data <= 32'h0011a700;
		52: data <= 32'h0014a702;
		53: data <= 32'h0018c140;
		54: data <= 32'h08000043;
		55: data <= 32'h0011a102;
		56: data <= 32'h0018c240;
		57: data <= 32'h08000043;
		58: data <= 32'h0315a020;
		59: data <= 32'hac540014;
		60: data <= 32'h200e0108;
		61: data <= 32'h200d0002;
		62: data <= 32'h016d5825;
		63: data <= 32'hac4b0008;
		64: data <= 32'h0018c202;
		65: data <= 32'h01c00008;
		66: data <= 32'h03400008;
		67: data <= 32'h1280001e;
		68: data <= 32'h2294ffff;
		69: data <= 32'h1280001e;
		70: data <= 32'h2294ffff;
		71: data <= 32'h1280001e;
		72: data <= 32'h2294ffff;
		73: data <= 32'h1280001e;
		74: data <= 32'h2294ffff;
		75: data <= 32'h1280001e;
		76: data <= 32'h2294ffff;
		77: data <= 32'h1280001e;
		78: data <= 32'h2294ffff;
		79: data <= 32'h1280001e;
		80: data <= 32'h2294ffff;
		81: data <= 32'h1280001e;
		82: data <= 32'h2294ffff;
		83: data <= 32'h1280001e;
		84: data <= 32'h2294ffff;
		85: data <= 32'h1280001e;
		86: data <= 32'h2294ffff;
		87: data <= 32'h1280001e;
		88: data <= 32'h2294ffff;
		89: data <= 32'h1280001e;
		90: data <= 32'h2294ffff;
		91: data <= 32'h1280001e;
		92: data <= 32'h2294ffff;
		93: data <= 32'h1280001e;
		94: data <= 32'h2294ffff;
		95: data <= 32'h1280001e;
		96: data <= 32'h2294ffff;
		97: data <= 32'h1280001e;
		98: data <= 32'h201500c0;
		99: data <= 32'h0800003a;
		100: data <= 32'h201500f9;
		101: data <= 32'h0800003a;
		102: data <= 32'h201500a4;
		103: data <= 32'h0800003a;
		104: data <= 32'h201500b0;
		105: data <= 32'h0800003a;
		106: data <= 32'h20150099;
		107: data <= 32'h0800003a;
		108: data <= 32'h20150092;
		109: data <= 32'h0800003a;
		110: data <= 32'h20150082;
		111: data <= 32'h0800003a;
		112: data <= 32'h201500f8;
		113: data <= 32'h0800003a;
		114: data <= 32'h20150080;
		115: data <= 32'h0800003a;
		116: data <= 32'h20150090;
		117: data <= 32'h0800003a;
		118: data <= 32'h20150088;
		119: data <= 32'h0800003a;
		120: data <= 32'h20150083;
		121: data <= 32'h0800003a;
		122: data <= 32'h201500c6;
		123: data <= 32'h0800003a;
		124: data <= 32'h201500a1;
		125: data <= 32'h0800003a;
		126: data <= 32'h20150086;
		127: data <= 32'h0800003a;
		128: data <= 32'h2015008e;
		129: data <= 32'h0800003a;
	endcase
endmodule
