`timescale 1ns/1ps

module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
	case(addr[10:2])	//Address Must Be Word Aligned.
0: data <= 32'b00001000000000000000000000000011;
1: data <= 32'b00001000000000000000000000100001;
2: data <= 32'b00001000000000000000000010000010;
3: data <= 32'b00100000000011100000000000100100;
4: data <= 32'b00111100000000100100000000000000;
5: data <= 32'b10101100010000000000000000001000;
6: data <= 32'b00100000000001001111110000011000;
7: data <= 32'b10101100010001000000000000000000;
8: data <= 32'b00000001110000000000000000001000;
9: data <= 32'b00100000000001001111111111111111;
10: data <= 32'b10101100010001000000000000000100;
11: data <= 32'b00100000000001010000000000000011;
12: data <= 32'b10101100010001010000000000001000;
13: data <= 32'b00100000000110000000000000001000;
14: data <= 32'b10001100010000110000000000011000;
15: data <= 32'b00100000011000111111111111111111;
16: data <= 32'b00011000011000001111111111111101;
17: data <= 32'b10001100010010000000000000011100;
18: data <= 32'b10001100010100000000000000011100;
19: data <= 32'b10001100010010010000000000100000;
20: data <= 32'b10001100010100010000000000100000;
21: data <= 32'b00000001000000000101000000100000;
22: data <= 32'b00000001010010010101000000100010;
23: data <= 32'b00011101010000001111111111111110;
24: data <= 32'b00010001010000000000000000000100;
25: data <= 32'b00000001010010010101000000100000;
26: data <= 32'b00000001001000000100000000100000;
27: data <= 32'b00000001010000000100100000100000;
28: data <= 32'b00001000000000000000000000010101;
29: data <= 32'b10101100010010010000000000100100;
30: data <= 32'b10101100010010010000000000001100;
31: data <= 32'b00000000100000000010000000100000;
32: data <= 32'b00001000000000000000000000011111;
33: data <= 32'b10001100010010110000000000001000;
34: data <= 32'b00110001011010111111111111111001;
35: data <= 32'b10101100010010110000000000001000;
36: data <= 32'b00100000000110010000000000001000;
37: data <= 32'b00010011000110010000000000001101;
38: data <= 32'b00000000000110011100100001000010;
39: data <= 32'b00010011000110010000000000001000;
40: data <= 32'b00000000000110011100100001000010;
41: data <= 32'b00010011000110010000000000000010;
42: data <= 32'b00000000000110011100100001000010;
43: data <= 32'b00010011000110010000000000001011;
44: data <= 32'b00000000000100001010011100000000;
45: data <= 32'b00000000000101001010011100000010;
46: data <= 32'b00000000000110001100001001000000;
47: data <= 32'b00001000000000000000000001000011;
48: data <= 32'b00000000000100001010000100000010;
49: data <= 32'b00000000000110001100001001000000;
50: data <= 32'b00001000000000000000000001000011;
51: data <= 32'b00000000000100011010011100000000;
52: data <= 32'b00000000000101001010011100000010;
53: data <= 32'b00000000000110001100000101000000;
54: data <= 32'b00001000000000000000000001000011;
55: data <= 32'b00000000000100011010000100000010;
56: data <= 32'b00000000000110001100001001000000;
57: data <= 32'b00001000000000000000000001000011;
58: data <= 32'b00000011000101011010000000100000;
59: data <= 32'b10101100010101000000000000010100;
60: data <= 32'b00100000000011100000000100001000;
61: data <= 32'b00100000000011010000000000000010;
62: data <= 32'b00000001011011010101100000100101;
63: data <= 32'b10101100010010110000000000001000;
64: data <= 32'b00000000000110001100001000000010;
65: data <= 32'b00000001110000000000000000001000;
66: data <= 32'b00000011010000000000000000001000;
67: data <= 32'b00010010100000000000000000011110;
68: data <= 32'b00100010100101001111111111111111;
69: data <= 32'b00010010100000000000000000011110;
70: data <= 32'b00100010100101001111111111111111;
71: data <= 32'b00010010100000000000000000011110;
72: data <= 32'b00100010100101001111111111111111;
73: data <= 32'b00010010100000000000000000011110;
74: data <= 32'b00100010100101001111111111111111;
75: data <= 32'b00010010100000000000000000011110;
76: data <= 32'b00100010100101001111111111111111;
77: data <= 32'b00010010100000000000000000011110;
78: data <= 32'b00100010100101001111111111111111;
79: data <= 32'b00010010100000000000000000011110;
80: data <= 32'b00100010100101001111111111111111;
81: data <= 32'b00010010100000000000000000011110;
82: data <= 32'b00100010100101001111111111111111;
83: data <= 32'b00010010100000000000000000011110;
84: data <= 32'b00100010100101001111111111111111;
85: data <= 32'b00010010100000000000000000011110;
86: data <= 32'b00100010100101001111111111111111;
87: data <= 32'b00010010100000000000000000011110;
88: data <= 32'b00100010100101001111111111111111;
89: data <= 32'b00010010100000000000000000011110;
90: data <= 32'b00100010100101001111111111111111;
91: data <= 32'b00010010100000000000000000011110;
92: data <= 32'b00100010100101001111111111111111;
93: data <= 32'b00010010100000000000000000011110;
94: data <= 32'b00100010100101001111111111111111;
95: data <= 32'b00010010100000000000000000011110;
96: data <= 32'b00100010100101001111111111111111;
97: data <= 32'b00010010100000000000000000011110;
98: data <= 32'b00100000000101010000000011000000;
99: data <= 32'b00001000000000000000000000111010;
100: data <= 32'b00100000000101010000000011111001;
101: data <= 32'b00001000000000000000000000111010;
102: data <= 32'b00100000000101010000000010100100;
103: data <= 32'b00001000000000000000000000111010;
104: data <= 32'b00100000000101010000000010110000;
105: data <= 32'b00001000000000000000000000111010;
106: data <= 32'b00100000000101010000000010011001;
107: data <= 32'b00001000000000000000000000111010;
108: data <= 32'b00100000000101010000000010010010;
109: data <= 32'b00001000000000000000000000111010;
110: data <= 32'b00100000000101010000000010000010;
111: data <= 32'b00001000000000000000000000111010;
112: data <= 32'b00100000000101010000000011111000;
113: data <= 32'b00001000000000000000000000111010;
114: data <= 32'b00100000000101010000000010000000;
115: data <= 32'b00001000000000000000000000111010;
116: data <= 32'b00100000000101010000000010010000;
117: data <= 32'b00001000000000000000000000111010;
118: data <= 32'b00100000000101010000000010001000;
119: data <= 32'b00001000000000000000000000111010;
120: data <= 32'b00100000000101010000000010000011;
121: data <= 32'b00001000000000000000000000111010;
122: data <= 32'b00100000000101010000000011000110;
123: data <= 32'b00001000000000000000000000111010;
124: data <= 32'b00100000000101010000000010100001;
125: data <= 32'b00001000000000000000000000111010;
126: data <= 32'b00100000000101010000000010000110;
127: data <= 32'b00001000000000000000000000111010;
128: data <= 32'b00100000000101010000000010001110;
129: data <= 32'b00001000000000000000000000111010;
130: data <= 32'b00000011010000000000000000001000;





		
	   default:	data <= 32'h0800_0000;
	endcase
endmodule
