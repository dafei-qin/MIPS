`timescale 1ns/1ps
module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];
always@(*)
	case(addr[10:2])
		0: data <= 32'h08000074;
		1: data <= 32'h08000003;
		2: data <= 32'h08000074;
		3: data <= 32'h3c014000;
		4: data <= 32'h20210008;
		5: data <= 32'hafa80004;
		6: data <= 32'hafa90008;
		7: data <= 32'hafaa000c;
		8: data <= 32'hafbf0010;
		9: data <= 32'h3c09ffff;
		10: data <= 32'h2529fff9;
		11: data <= 32'h8c280000;
		12: data <= 32'h01094024;
		13: data <= 32'hac280000;
		14: data <= 32'h3c010000;
		15: data <= 32'h24210400;
		16: data <= 32'h8c28fffc;
		17: data <= 32'h3c014000;
		18: data <= 32'h20210014;
		19: data <= 32'h2409000f;
		20: data <= 32'h01284824;
		21: data <= 32'h0c000035;
		22: data <= 32'h21290100;
		23: data <= 32'hac290000;
		24: data <= 32'h240900f0;
		25: data <= 32'h01284824;
		26: data <= 32'h00094902;
		27: data <= 32'h0c000035;
		28: data <= 32'h21290200;
		29: data <= 32'hac290000;
		30: data <= 32'h24090f00;
		31: data <= 32'h01284824;
		32: data <= 32'h00094a02;
		33: data <= 32'h0c000035;
		34: data <= 32'h21290400;
		35: data <= 32'hac290000;
		36: data <= 32'h2409f000;
		37: data <= 32'h01284824;
		38: data <= 32'h00094b02;
		39: data <= 32'h0c000035;
		40: data <= 32'h21290800;
		41: data <= 32'hac290000;
		42: data <= 32'h3c014000;
		43: data <= 32'h20210008;
		44: data <= 32'h8c290000;
		45: data <= 32'h200a0002;
		46: data <= 32'h012a4825;
		47: data <= 32'hac290000;
		48: data <= 32'h8fa80004;
		49: data <= 32'h8fa90008;
		50: data <= 32'h8faa000c;
		51: data <= 32'h8fbf0010;
		52: data <= 32'h03400008;
		53: data <= 32'h1120001e;
		54: data <= 32'h2129ffff;
		55: data <= 32'h1120001e;
		56: data <= 32'h2129ffff;
		57: data <= 32'h1120001e;
		58: data <= 32'h2129ffff;
		59: data <= 32'h1120001e;
		60: data <= 32'h2129ffff;
		61: data <= 32'h1120001e;
		62: data <= 32'h2129ffff;
		63: data <= 32'h1120001e;
		64: data <= 32'h2129ffff;
		65: data <= 32'h1120001e;
		66: data <= 32'h2129ffff;
		67: data <= 32'h1120001e;
		68: data <= 32'h2129ffff;
		69: data <= 32'h1120001e;
		70: data <= 32'h2129ffff;
		71: data <= 32'h1120001e;
		72: data <= 32'h2129ffff;
		73: data <= 32'h1120001e;
		74: data <= 32'h2129ffff;
		75: data <= 32'h1120001e;
		76: data <= 32'h2129ffff;
		77: data <= 32'h1120001e;
		78: data <= 32'h2129ffff;
		79: data <= 32'h1120001e;
		80: data <= 32'h2129ffff;
		81: data <= 32'h1120001e;
		82: data <= 32'h2129ffff;
		83: data <= 32'h1120001e;
		84: data <= 32'h240900c0;
		85: data <= 32'h03e00008;
		86: data <= 32'h240900f9;
		87: data <= 32'h03e00008;
		88: data <= 32'h240900a4;
		89: data <= 32'h03e00008;
		90: data <= 32'h240900b0;
		91: data <= 32'h03e00008;
		92: data <= 32'h24090099;
		93: data <= 32'h03e00008;
		94: data <= 32'h24090092;
		95: data <= 32'h03e00008;
		96: data <= 32'h24090082;
		97: data <= 32'h03e00008;
		98: data <= 32'h240900f8;
		99: data <= 32'h03e00008;
		100: data <= 32'h24090080;
		101: data <= 32'h03e00008;
		102: data <= 32'h24090090;
		103: data <= 32'h03e00008;
		104: data <= 32'h24090088;
		105: data <= 32'h03e00008;
		106: data <= 32'h24090083;
		107: data <= 32'h03e00008;
		108: data <= 32'h240900c6;
		109: data <= 32'h03e00008;
		110: data <= 32'h240900a1;
		111: data <= 32'h03e00008;
		112: data <= 32'h24090086;
		113: data <= 32'h03e00008;
		114: data <= 32'h2409008e;
		115: data <= 32'h03e00008;
		116: data <= 32'hafa80004;
		117: data <= 32'h3c084000;
		118: data <= 32'h21080010;
		119: data <= 32'h8d010000;
		120: data <= 32'h3c084000;
		121: data <= 32'h2108000c;
		122: data <= 32'h10200003;
		123: data <= 32'h20010001;
		124: data <= 32'had010000;
		125: data <= 32'h08000080;
		126: data <= 32'h20010000;
		127: data <= 32'had010000;
		128: data <= 32'h8fa80004;
		129: data <= 32'h20010002;
		130: data <= 32'hafa80004;
		131: data <= 32'h3c084000;
		132: data <= 32'h21080020;
		133: data <= 32'had010000;
		134: data <= 32'h8d010000;
		135: data <= 32'h2021fff6;
		136: data <= 32'h1420fffd;
		137: data <= 32'h8d05fffc;
		138: data <= 32'h20010000;
		139: data <= 32'had010000;
		140: data <= 32'h8fa80004;
		141: data <= 32'hafa80004;
		142: data <= 32'h3c084000;
		143: data <= 32'h21080010;
		144: data <= 32'h8d010000;
		145: data <= 32'h3c084000;
		146: data <= 32'h2108000c;
		147: data <= 32'h10200003;
		148: data <= 32'h20010000;
		149: data <= 32'had010000;
		150: data <= 32'h08000099;
		151: data <= 32'h20010000;
		152: data <= 32'had010000;
		153: data <= 32'h8fa80004;
		154: data <= 32'hafa80004;
		155: data <= 32'h3c084000;
		156: data <= 32'h21080010;
		157: data <= 32'h8d010000;
		158: data <= 32'h3c084000;
		159: data <= 32'h2108000c;
		160: data <= 32'h10200003;
		161: data <= 32'h20010001;
		162: data <= 32'had010000;
		163: data <= 32'h080000a6;
		164: data <= 32'h20010000;
		165: data <= 32'had010000;
		166: data <= 32'h8fa80004;
		167: data <= 32'h20010002;
		168: data <= 32'hafa80004;
		169: data <= 32'h3c084000;
		170: data <= 32'h21080020;
		171: data <= 32'had010000;
		172: data <= 32'h8d010000;
		173: data <= 32'h2021fff6;
		174: data <= 32'h1420fffd;
		175: data <= 32'h8d06fffc;
		176: data <= 32'h20010000;
		177: data <= 32'had010000;
		178: data <= 32'h8fa80004;
		179: data <= 32'hafa80004;
		180: data <= 32'h3c084000;
		181: data <= 32'h21080010;
		182: data <= 32'h8d010000;
		183: data <= 32'h3c084000;
		184: data <= 32'h2108000c;
		185: data <= 32'h10200003;
		186: data <= 32'h20010000;
		187: data <= 32'had010000;
		188: data <= 32'h080000bf;
		189: data <= 32'h20010000;
		190: data <= 32'had010000;
		191: data <= 32'h8fa80004;
		192: data <= 32'h3c014000;
		193: data <= 32'h20210008;
		194: data <= 32'hac200000;
		195: data <= 32'hafa80004;
		196: data <= 32'hafa90008;
		197: data <= 32'h3c010000;
		198: data <= 32'h24210400;
		199: data <= 32'h3c09ff00;
		200: data <= 32'h00094c02;
		201: data <= 32'h8c28fffc;
		202: data <= 32'h01094024;
		203: data <= 32'h01054020;
		204: data <= 32'hac28fffc;
		205: data <= 32'h3c014000;
		206: data <= 32'h20210008;
		207: data <= 32'h2408d8ef;
		208: data <= 32'hac28fff8;
		209: data <= 32'hac28fffc;
		210: data <= 32'h20080003;
		211: data <= 32'hac280000;
		212: data <= 32'h8fa80004;
		213: data <= 32'h8fa90008;
		214: data <= 32'h3c014000;
		215: data <= 32'h20210008;
		216: data <= 32'hac200000;
		217: data <= 32'hafa80004;
		218: data <= 32'hafa90008;
		219: data <= 32'h3c010000;
		220: data <= 32'h24210400;
		221: data <= 32'h3c0800ff;
		222: data <= 32'h00084402;
		223: data <= 32'h3c09ffff;
		224: data <= 32'h01284820;
		225: data <= 32'h8c28fffc;
		226: data <= 32'h00063200;
		227: data <= 32'h01284024;
		228: data <= 32'h01064020;
		229: data <= 32'h00063202;
		230: data <= 32'hac28fffc;
		231: data <= 32'h3c014000;
		232: data <= 32'h20210008;
		233: data <= 32'h2008d8ef;
		234: data <= 32'hac28fff8;
		235: data <= 32'hac28fffc;
		236: data <= 32'h20080003;
		237: data <= 32'hac280000;
		238: data <= 32'h8fa80004;
		239: data <= 32'h8fa90008;
		240: data <= 32'h00c55820;
		241: data <= 32'hafa80004;
		242: data <= 32'h3c084000;
		243: data <= 32'h21080010;
		244: data <= 32'h8d010000;
		245: data <= 32'h3c084000;
		246: data <= 32'h2108000c;
		247: data <= 32'h10200003;
		248: data <= 32'h20010002;
		249: data <= 32'had010000;
		250: data <= 32'h080000fd;
		251: data <= 32'h20010000;
		252: data <= 32'had010000;
		253: data <= 32'h8fa80004;
		254: data <= 32'hafa80004;
		255: data <= 32'h3c084000;
		256: data <= 32'h21080020;
		257: data <= 32'h8d010000;
		258: data <= 32'h1420fffe;
		259: data <= 32'had0bfff8;
		260: data <= 32'h20010001;
		261: data <= 32'had010000;
		262: data <= 32'h8d010000;
		263: data <= 32'h2021ffeb;
		264: data <= 32'h1420fffd;
		265: data <= 32'had000000;
		266: data <= 32'h8fa80004;
		267: data <= 32'hafa80004;
		268: data <= 32'h3c084000;
		269: data <= 32'h21080010;
		270: data <= 32'h8d010000;
		271: data <= 32'h3c084000;
		272: data <= 32'h2108000c;
		273: data <= 32'h10200003;
		274: data <= 32'h20010000;
		275: data <= 32'had010000;
		276: data <= 32'h08000117;
		277: data <= 32'h20010000;
		278: data <= 32'had010000;
		279: data <= 32'h8fa80004;
		280: data <= 32'h08000118;
	endcase
endmodule
