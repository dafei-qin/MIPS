`timescale 1ns/1ps
module ALU_tb;
reg [31:0] A, B;
reg [5:0] ALUFun;
reg Sign;
wire [31:0] Z;
ALU test(A, B, ALUFun, Sign, Z, S, V);

initial begin
/*
	Sign = 1;
	A = 32'b10000000000000000000000000000000;
	B = 32'b10000000000000000000000000000000;
	ALUFun = 6'b110011;
	#1
	ALUFun = 6'b110001;
	#1
	A = 32'b10000000000000000000000000000000;
	B = 32'b01111111111111111111111111111111;
	ALUFun = 6'b110101;
	#1
	A = 32'b00000000000000000000000000000000;
	B = 32'b00000000000000000000000000000000;
	ALUFun = 6'b111101;
	#1
	ALUFun = 6'b111011;
	#1
	ALUFun = 6'b111111;
*/
	A = 32'b10000000000000000000000000011101;
	B = 32'b10000000000000000000000000000001;
	ALUFun = 6'b100000;
	#1
	A = 32'b1000000000000000000000000000011;
	ALUFun = 6'b100001;
	#1
	ALUFun = 6'b100011;
end

endmodule